`timescale 1ns / 1ps

module digital_stopwatchtb(

    );
endmodule
